module mymodule(input A1, input A2, output [7:0] cout);
    input A1, A2;
    reg cout;

    

endmodule

